module bin_2_bcd (carryout,out,d,u);
  input carryout;
  input [3:0] out;
  output [1:0]d;
  output [3:0]u;
  wire s0;
  wire s1;
  wire s2;
  wire s3;
  assign d[1] = ((carryout & out[2]) | (carryout & out[3]));
  assign s0 = ~ carryout;
  assign s1 = ~ out[3];
  assign s2 = ~ out[2];
  assign s3 = ~ out[1];
  assign d[0] = ((s0 & out[3] & out[1]) | (s0 & out[3] & out[2]) | (carryout & s1 & s2) | (out[3] & out[1] & out[2]));
  assign u[3] = ((s0 & out[3] & s3 & s2) | (carryout & s1 & out[1] & s2) | (carryout & out[3] & s3 & out[2]));
  assign u[2] = ((s0 & s1 & out[2]) | (s0 & out[1] & out[2]) | (carryout & s3 & s2) | (carryout & out[3] & s2));
  assign u[1] = ((carryout & out[0] & out[1] & out[2]) | (s0 & out[3] & s3 & out[2]) | (carryout & s1 & s3 & s2) | (carryout & out[3] & out[1] & s2) | (s0 & s1 & out[1]) | (s1 & out[1] & out[2]));
  assign u[0] = ((s0 & out[0]) | (s1 & out[0]) | (out[0] & s3) | (out[0] & s2));
endmodule
